CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 1520 1 120 10
176 79 1364 717
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 175 457 272
9437202 0
0
6 Title:
5 Name:
0
0
0
59
13 Logic Switch~
5 123 1186 0 10 11
0 25 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V8
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7100 0 0
2
41141.7 1
0
13 Logic Switch~
5 175 780 0 10 11
0 32 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3820 0 0
2
41141.6 0
0
13 Logic Switch~
5 180 329 0 10 11
0 36 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7678 0 0
2
41141.6 0
0
12 Hex Display~
7 394 1640 0 18 19
10 5 4 2 6 0 0 0 0 0
0 1 0 1 1 0 1 1 5
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP3
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
961 0 0
2
41141.7 11
0
14 Logic Display~
6 576 1695 0 1 2
10 6
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L20
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3178 0 0
2
41141.7 10
0
14 Logic Display~
6 470 1701 0 1 2
10 2
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L19
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3409 0 0
2
41141.7 9
0
14 Logic Display~
6 360 1706 0 1 2
10 4
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L18
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3951 0 0
2
41141.7 8
0
14 Logic Display~
6 253 1713 0 1 2
10 5
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L17
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8885 0 0
2
41141.7 7
0
2 +V
167 128 1764 0 1 3
0 8
0
0 0 54256 0
3 10V
-11 -22 10 -14
3 V12
-10 -32 11 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
3780 0 0
2
41141.7 6
0
6 JK RN~
219 533 1821 0 6 22
0 8 2 8 3 43 6
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
4 U12B
-14 -42 14 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 512 2 2 12 0
1 U
9265 0 0
2
41141.7 5
0
6 JK RN~
219 425 1830 0 6 22
0 8 4 8 3 44 2
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
4 U12A
-14 -42 14 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 512 2 1 12 0
1 U
9442 0 0
2
41141.7 4
0
6 JK RN~
219 318 1839 0 6 22
0 8 5 8 3 45 4
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
4 U11B
-14 -42 14 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 512 2 2 11 0
1 U
9424 0 0
2
41141.7 3
0
6 JK RN~
219 218 1848 0 6 22
0 8 7 8 3 46 5
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
4 U11A
-14 -42 14 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 512 2 1 11 0
1 U
9968 0 0
2
41141.7 2
0
10 2-In NAND~
219 245 1925 0 3 22
0 4 2 3
0
0 0 624 512
4 7400
-7 -24 21 -16
4 U10B
-11 -25 17 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 10 0
1 U
9281 0 0
2
41141.7 1
0
7 Pulser~
4 140 1840 0 10 12
0 47 48 49 7 0 0 5 5 5
8
0
0 0 4656 0
0
3 V10
-10 -28 11 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
8464 0 0
2
41141.7 0
0
7 Pulser~
4 168 252 0 10 12
0 50 51 52 41 0 0 5 5 5
8
0
0 0 4656 0
0
2 V2
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
7168 0 0
2
41141.7 0
0
7 Pulser~
4 138 703 0 10 12
0 53 54 55 34 0 0 5 5 5
8
0
0 0 4656 0
0
2 V5
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
3171 0 0
2
41141.7 0
0
7 Pulser~
4 165 1467 0 10 12
0 56 57 58 14 0 0 5 5 5
8
0
0 0 4656 0
0
2 V9
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
4139 0 0
2
41141.7 0
0
10 2-In NAND~
219 270 1552 0 3 22
0 11 10 9
0
0 0 624 512
4 7400
-7 -24 21 -16
4 U10A
-11 -25 17 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 10 0
1 U
6435 0 0
2
41141.7 0
0
6 JK RN~
219 243 1475 0 6 22
0 15 14 15 9 59 12
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U9B
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 512 2 2 9 0
1 U
5283 0 0
2
41141.7 11
0
6 JK RN~
219 343 1466 0 6 22
0 15 12 15 9 60 11
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U9A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 512 2 1 9 0
1 U
6874 0 0
2
41141.7 10
0
6 JK RN~
219 450 1457 0 6 22
0 15 11 15 9 61 13
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U8B
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 512 2 2 8 0
1 U
5305 0 0
2
41141.7 9
0
6 JK RN~
219 558 1448 0 6 22
0 15 13 15 9 62 10
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U8A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 512 2 1 8 0
1 U
34 0 0
2
41141.7 8
0
2 +V
167 153 1391 0 1 3
0 15
0
0 0 54256 0
3 10V
-11 -22 10 -14
3 V11
-10 -32 11 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
969 0 0
2
41141.7 7
0
14 Logic Display~
6 278 1340 0 1 2
10 12
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L16
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8402 0 0
2
41141.7 6
0
14 Logic Display~
6 385 1333 0 1 2
10 11
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L15
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3751 0 0
2
41141.7 5
0
14 Logic Display~
6 495 1328 0 1 2
10 13
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L14
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4292 0 0
2
41141.7 4
0
14 Logic Display~
6 601 1322 0 1 2
10 10
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L13
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6118 0 0
2
41141.7 3
0
12 Hex Display~
7 419 1267 0 18 19
10 12 11 13 10 0 0 0 0 0
0 1 1 1 0 0 0 0 7
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP4
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
34 0 0
2
41141.7 2
0
7 Pulser~
4 96 1105 0 10 12
0 63 64 65 20 0 0 5 5 5
8
0
0 0 4656 0
0
2 V7
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
6357 0 0
2
41141.7 0
0
9 Inverter~
13 184 1083 0 2 22
0 16 24
0
0 0 624 270
6 74LS04
-21 -19 21 -11
3 U7A
16 -8 37 0
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 7 0
1 U
319 0 0
2
41141.7 0
0
14 Logic Display~
6 424 973 0 1 2
10 16
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L12
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3976 0 0
2
41141.7 10
0
14 Logic Display~
6 410 973 0 1 2
10 17
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L11
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7634 0 0
2
41141.7 9
0
14 Logic Display~
6 395 973 0 1 2
10 18
0
0 0 53872 0
6 100MEG
3 -16 45 -8
3 L10
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
523 0 0
2
41141.7 8
0
14 Logic Display~
6 381 973 0 1 2
10 19
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L9
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6748 0 0
2
41141.7 7
0
6 JK RN~
219 562 1115 0 6 22
0 17 20 21 25 66 16
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U6B
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 512 2 2 6 0
1 U
6901 0 0
2
41141.7 5
0
6 JK RN~
219 461 1115 0 6 22
0 18 20 22 25 21 17
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U6A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 0 2 1 6 0
1 U
842 0 0
2
41141.7 4
0
6 JK RN~
219 353 1115 0 6 22
0 19 20 23 25 22 18
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U5B
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 0 2 2 5 0
1 U
3277 0 0
2
41141.7 3
0
6 JK RN~
219 261 1115 0 6 22
0 16 20 24 25 23 19
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U5A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 0 2 1 5 0
1 U
4212 0 0
2
41141.7 2
0
6 JK RN~
219 261 711 0 6 22
0 35 34 35 32 31 27
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U4B
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 0 2 2 4 0
1 U
4720 0 0
2
41141.6 11
0
6 JK RN~
219 361 702 0 6 22
0 35 31 35 32 30 33
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U4A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 0 2 1 4 0
1 U
5551 0 0
2
41141.6 10
0
6 JK RN~
219 469 694 0 6 22
0 35 30 35 32 29 28
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U3B
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 0 2 2 3 0
1 U
6986 0 0
2
41141.6 9
0
6 JK RN~
219 567 684 0 6 22
0 35 29 35 32 67 26
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U3A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 512 2 1 3 0
1 U
8745 0 0
2
41141.6 8
0
2 +V
167 171 627 0 1 3
0 35
0
0 0 54256 0
3 10V
-11 -22 10 -14
2 V6
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
9592 0 0
2
41141.6 7
0
14 Logic Display~
6 296 576 0 1 2
10 27
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
8748 0 0
2
41141.6 6
0
14 Logic Display~
6 403 569 0 1 2
10 33
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
7168 0 0
2
41141.6 5
0
14 Logic Display~
6 513 563 0 1 2
10 28
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
631 0 0
2
41141.6 4
0
14 Logic Display~
6 619 558 0 1 2
10 26
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9466 0 0
2
41141.6 3
0
12 Hex Display~
7 437 486 0 18 19
10 27 33 28 26 0 0 0 0 0
0 0 1 1 0 0 0 0 1
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP2
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
3266 0 0
2
41141.6 2
0
12 Hex Display~
7 442 52 0 18 19
10 37 38 39 40 0 0 0 0 0
0 1 0 0 0 1 1 1 15
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
7693 0 0
2
41141.6 0
0
14 Logic Display~
6 624 107 0 1 2
10 40
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3723 0 0
2
41141.6 0
0
14 Logic Display~
6 518 113 0 1 2
10 39
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3440 0 0
2
41141.6 0
0
14 Logic Display~
6 408 118 0 1 2
10 38
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
6263 0 0
2
41141.6 0
0
14 Logic Display~
6 301 125 0 1 2
10 37
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4900 0 0
2
41141.6 0
0
2 +V
167 176 176 0 1 3
0 42
0
0 0 54256 0
3 10V
-11 -22 10 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
8783 0 0
2
41141.6 0
0
6 JK RN~
219 581 233 0 6 22
0 42 39 42 36 68 40
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U2B
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 512 2 2 2 0
1 U
3221 0 0
2
41141.6 0
0
6 JK RN~
219 473 242 0 6 22
0 42 38 42 36 69 39
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U2A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 512 2 1 2 0
1 U
3215 0 0
2
41141.6 0
0
6 JK RN~
219 366 251 0 6 22
0 42 37 42 36 70 38
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U1B
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 512 2 2 1 0
1 U
7903 0 0
2
41141.6 0
0
6 JK RN~
219 266 260 0 6 22
0 42 41 42 36 71 37
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U1A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 512 2 1 1 0
1 U
7121 0 0
2
41141.6 0
0
121
0 2 2 0 0 12432 0 0 14 12 0 4
470 1813
471 1813
471 1934
271 1934
4 0 3 0 0 0 0 13 0 0 3 2
218 1879
218 1879
4 3 3 0 0 8320 0 10 14 0 0 7
533 1852
533 1898
218 1898
218 1879
218 1879
218 1925
220 1925
0 1 4 0 0 4096 0 0 14 13 0 3
360 1822
360 1916
271 1916
4 0 3 0 0 0 0 11 0 0 3 2
425 1861
425 1898
4 0 3 0 0 0 0 12 0 0 3 2
318 1870
318 1898
1 0 5 0 0 8320 0 4 0 0 14 3
403 1664
403 1751
253 1751
2 0 4 0 0 0 0 4 0 0 13 3
397 1664
397 1744
360 1744
3 0 2 0 0 0 0 4 0 0 12 3
391 1664
391 1737
470 1737
4 0 6 0 0 8320 0 4 0 0 11 3
385 1664
385 1730
598 1730
1 6 6 0 0 0 0 5 10 0 0 4
576 1713
598 1713
598 1804
557 1804
1 0 2 0 0 0 0 6 0 0 24 2
470 1719
470 1813
1 0 4 0 0 4224 0 7 0 0 25 2
360 1724
360 1822
0 1 5 0 0 0 0 0 8 26 0 2
253 1831
253 1731
4 2 7 0 0 4224 0 15 13 0 0 2
170 1840
187 1840
1 0 8 0 0 4096 0 13 0 0 17 4
194 1831
181 1831
181 1832
176 1832
3 0 8 0 0 8192 0 13 0 0 23 3
194 1849
176 1849
176 1773
1 0 8 0 0 0 0 12 0 0 19 2
294 1822
274 1822
3 0 8 0 0 0 0 12 0 0 23 3
294 1840
274 1840
274 1773
1 0 8 0 0 0 0 11 0 0 21 4
401 1813
384 1813
384 1814
387 1814
3 0 8 0 0 0 0 11 0 0 23 3
401 1831
387 1831
387 1773
1 0 8 0 0 0 0 10 0 0 23 2
509 1804
493 1804
1 3 8 0 0 4224 0 9 10 0 0 4
128 1773
493 1773
493 1822
509 1822
6 2 2 0 0 0 0 11 10 0 0 2
449 1813
502 1813
6 2 4 0 0 0 0 12 11 0 0 2
342 1822
394 1822
6 2 5 0 0 0 0 13 12 0 0 2
242 1831
287 1831
4 0 9 0 0 0 0 20 0 0 28 2
243 1506
243 1506
4 3 9 0 0 8320 0 23 19 0 0 7
558 1479
558 1525
243 1525
243 1506
243 1506
243 1552
245 1552
0 2 10 0 0 12416 0 0 19 37 0 4
601 1431
602 1431
602 1561
296 1561
0 1 11 0 0 4096 0 0 19 39 0 3
385 1449
385 1543
296 1543
4 0 9 0 0 0 0 22 0 0 28 2
450 1488
450 1525
4 0 9 0 0 0 0 21 0 0 28 2
343 1497
343 1525
1 0 12 0 0 8320 0 29 0 0 40 3
428 1291
428 1378
278 1378
2 0 11 0 0 0 0 29 0 0 39 3
422 1291
422 1371
385 1371
3 0 13 0 0 8192 0 29 0 0 38 3
416 1291
416 1364
495 1364
4 0 10 0 0 0 0 29 0 0 37 3
410 1291
410 1357
601 1357
1 6 10 0 0 0 0 28 23 0 0 3
601 1340
601 1431
582 1431
1 0 13 0 0 4224 0 27 0 0 50 2
495 1346
495 1440
1 0 11 0 0 4224 0 26 0 0 51 2
385 1351
385 1449
0 1 12 0 0 0 0 0 25 52 0 2
278 1458
278 1358
4 2 14 0 0 4224 0 18 20 0 0 2
195 1467
212 1467
1 0 15 0 0 4096 0 20 0 0 43 4
219 1458
206 1458
206 1459
201 1459
3 0 15 0 0 8192 0 20 0 0 49 3
219 1476
201 1476
201 1400
1 0 15 0 0 0 0 21 0 0 45 2
319 1449
299 1449
3 0 15 0 0 0 0 21 0 0 49 3
319 1467
299 1467
299 1400
1 0 15 0 0 0 0 22 0 0 47 4
426 1440
409 1440
409 1441
412 1441
3 0 15 0 0 0 0 22 0 0 49 3
426 1458
412 1458
412 1400
1 0 15 0 0 0 0 23 0 0 49 2
534 1431
518 1431
1 3 15 0 0 4224 0 24 23 0 0 4
153 1400
518 1400
518 1449
534 1449
6 2 13 0 0 0 0 22 23 0 0 2
474 1440
527 1440
6 2 11 0 0 0 0 21 22 0 0 2
367 1449
419 1449
6 2 12 0 0 0 0 20 21 0 0 2
267 1458
312 1458
0 0 16 0 0 8320 0 0 0 68 60 3
201 1048
201 1031
612 1031
1 0 17 0 0 8320 0 33 0 0 62 4
410 991
410 1083
507 1083
507 1098
1 0 18 0 0 4224 0 34 0 0 64 4
395 991
395 1083
397 1083
397 1098
1 0 19 0 0 4224 0 35 0 0 66 4
381 991
381 1083
304 1083
304 1098
2 0 20 0 0 8192 0 38 0 0 59 3
322 1107
305 1107
305 1161
2 0 20 0 0 0 0 37 0 0 59 3
430 1107
411 1107
411 1161
0 2 20 0 0 8320 0 0 36 73 0 5
174 1107
174 1161
514 1161
514 1107
531 1107
6 1 16 0 0 128 0 36 32 0 0 5
586 1098
612 1098
612 1031
424 1031
424 991
5 3 21 0 0 4224 0 37 36 0 0 2
491 1116
538 1116
6 1 17 0 0 128 0 37 36 0 0 2
485 1098
538 1098
5 3 22 0 0 4224 0 38 37 0 0 2
383 1116
437 1116
6 1 18 0 0 128 0 38 37 0 0 2
377 1098
437 1098
3 5 23 0 0 4224 0 38 39 0 0 2
329 1116
291 1116
6 1 19 0 0 128 0 39 38 0 0 2
285 1098
329 1098
2 3 24 0 0 8320 0 31 39 0 0 3
187 1101
187 1116
237 1116
1 1 16 0 0 128 0 39 31 0 0 5
237 1098
215 1098
215 1048
187 1048
187 1065
4 0 25 0 0 4096 0 37 0 0 72 2
461 1146
461 1185
4 0 25 0 0 0 0 38 0 0 72 4
353 1146
353 1170
354 1170
354 1185
4 0 25 0 0 0 0 39 0 0 72 2
261 1146
261 1185
4 1 25 0 0 8320 0 36 1 0 0 5
562 1146
562 1185
261 1185
261 1186
135 1186
4 2 20 0 0 128 0 30 39 0 0 4
126 1105
174 1105
174 1107
230 1107
1 6 26 0 0 8192 0 48 43 0 0 4
619 576
623 576
623 667
591 667
6 1 27 0 0 8192 0 40 45 0 0 3
285 694
296 694
296 594
1 6 28 0 0 8320 0 47 42 0 0 4
513 581
504 581
504 677
493 677
5 2 29 0 0 4224 0 42 43 0 0 4
499 695
519 695
519 676
536 676
5 2 30 0 0 12416 0 41 42 0 0 4
391 703
412 703
412 686
438 686
5 2 31 0 0 12416 0 40 41 0 0 4
291 712
305 712
305 694
330 694
4 0 32 0 0 4096 0 42 0 0 88 4
469 725
469 765
468 765
468 780
4 0 32 0 0 4096 0 41 0 0 88 2
361 733
361 780
4 0 32 0 0 0 0 40 0 0 88 4
261 742
261 765
262 765
262 780
1 0 27 0 0 8320 0 49 0 0 75 3
446 510
446 614
296 614
2 0 33 0 0 4096 0 49 0 0 87 3
440 510
440 607
395 607
3 0 28 0 0 0 0 49 0 0 76 3
434 510
434 600
504 600
4 0 26 0 0 8320 0 49 0 0 74 3
428 510
428 593
623 593
1 6 33 0 0 8320 0 46 41 0 0 4
403 587
395 587
395 685
385 685
4 1 32 0 0 8320 0 43 2 0 0 3
567 715
567 780
187 780
4 2 34 0 0 4224 0 17 40 0 0 2
168 703
230 703
1 0 35 0 0 4096 0 40 0 0 91 2
237 694
219 694
3 0 35 0 0 8192 0 40 0 0 97 3
237 712
219 712
219 636
1 0 35 0 0 0 0 41 0 0 93 2
337 685
317 685
3 0 35 0 0 0 0 41 0 0 97 3
337 703
317 703
317 636
1 0 35 0 0 0 0 42 0 0 95 4
445 677
437 677
437 676
430 676
3 0 35 0 0 0 0 42 0 0 97 3
445 695
430 695
430 636
1 0 35 0 0 0 0 43 0 0 97 2
543 667
525 667
1 3 35 0 0 4224 0 44 43 0 0 4
171 636
525 636
525 685
543 685
4 0 36 0 0 4096 0 57 0 0 109 2
473 273
473 329
4 0 36 0 0 0 0 58 0 0 109 2
366 282
366 329
4 0 36 0 0 0 0 59 0 0 109 4
266 291
266 324
267 324
267 329
1 0 37 0 0 8320 0 50 0 0 108 3
451 76
451 163
301 163
2 0 38 0 0 4096 0 50 0 0 107 3
445 76
445 156
408 156
3 0 39 0 0 8192 0 50 0 0 106 3
439 76
439 149
518 149
4 0 40 0 0 8320 0 50 0 0 105 3
433 76
433 142
624 142
1 6 40 0 0 0 0 51 56 0 0 3
624 125
624 216
605 216
1 0 39 0 0 4224 0 52 0 0 119 2
518 131
518 225
1 0 38 0 0 4224 0 53 0 0 120 2
408 136
408 234
0 1 37 0 0 0 0 0 54 121 0 2
301 243
301 143
4 1 36 0 0 8320 0 56 3 0 0 3
581 264
581 329
192 329
4 2 41 0 0 4224 0 16 59 0 0 2
198 252
235 252
1 0 42 0 0 4096 0 59 0 0 112 4
242 243
229 243
229 244
224 244
3 0 42 0 0 8192 0 59 0 0 118 3
242 261
224 261
224 185
1 0 42 0 0 0 0 58 0 0 114 2
342 234
322 234
3 0 42 0 0 0 0 58 0 0 118 3
342 252
322 252
322 185
1 0 42 0 0 0 0 57 0 0 116 4
449 225
432 225
432 226
435 226
3 0 42 0 0 0 0 57 0 0 118 3
449 243
435 243
435 185
1 0 42 0 0 0 0 56 0 0 118 2
557 216
541 216
1 3 42 0 0 4224 0 55 56 0 0 4
176 185
541 185
541 234
557 234
6 2 39 0 0 0 0 57 56 0 0 2
497 225
550 225
6 2 38 0 0 0 0 58 57 0 0 2
390 234
442 234
6 2 37 0 0 0 0 59 58 0 0 2
290 243
335 243
8
-32 0 0 0 700 0 0 0 0 3 2 1 2
3 LCD
0 0 0 7
244 1632 367 1673
249 1637 361 1668
7 Counter
-32 0 0 0 700 0 0 0 0 3 2 1 2
3 LCD
0 0 0 4
96 1632 176 1676
102 1639 169 1671
4 Mode
-96 0 0 0 700 255 0 0 0 3 2 1 2
3 LCD
0 0 0 2
129 1596 242 1725
136 1603 234 1698
2 10
-96 0 0 0 700 255 0 0 0 3 2 1 2
3 LCD
0 0 0 2
154 1223 267 1352
161 1230 259 1325
2 10
-32 0 0 0 700 0 0 0 0 3 2 1 2
3 LCD
0 0 0 4
121 1259 201 1303
127 1266 194 1298
4 Mode
-32 0 0 0 700 0 0 0 0 3 2 1 2
3 LCD
0 0 0 7
269 1259 392 1300
274 1264 386 1295
7 Counter
-32 0 0 0 700 0 0 0 0 3 2 1 2
3 LCD
0 0 0 7
260 45 383 86
265 50 377 81
7 Counter
-32 0 0 0 700 0 0 0 0 3 2 1 2
3 LCD
0 0 0 10
201 493 367 534
208 498 359 529
10 Count Down
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 1e-06 1e-07 1e-07
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
14112 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
