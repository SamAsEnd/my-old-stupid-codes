CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
90 0 30 90 10
94 79 1302 747
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
262 175 375 272
9437202 0
0
6 Title:
5 Name:
0
0
0
24
13 Logic Switch~
5 147 275 0 10 11
0 5 0 0 0 0 0 0 0 0
1
0
0 0 29424 0
2 5V
-6 -16 8 -8
1 A
-3 -26 4 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5130 0 0
2
41149 0
0
12 Hex Display~
7 501 146 0 16 19
10 2 4 22 23 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
2 D4
-8 -38 6 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 512 0 0 0 0
4 DISP
391 0 0
2
41149.1 0
0
9 2-In AND~
219 889 406 0 3 22
0 7 6 8
0
0 0 624 90
6 74LS08
-21 -24 21 -16
2 AD
19 -5 33 3
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 7 0
1 U
3124 0 0
2
41149.1 0
0
10 2-In NAND~
219 962 501 0 3 22
0 4 3 7
0
0 0 624 512
4 7400
-7 -24 21 -16
3 ND4
-8 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
3421 0 0
2
41149.1 0
0
6 JK RN~
219 1266 339 0 6 22
0 5 9 5 7 24 2
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
4 JK12
-14 -42 14 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 512 2 2 17 0
1 U
8157 0 0
2
41149.1 1
0
6 JK RN~
219 1344 339 0 6 22
0 5 2 5 7 25 4
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
4 JK13
-14 -42 14 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 512 2 1 19 0
1 U
5572 0 0
2
41149.1 0
0
10 2-In NAND~
219 961 436 0 3 22
0 10 9 6
0
0 0 624 512
4 7400
-7 -24 21 -16
3 ND3
-8 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 0 0
1 U
8901 0 0
2
41149.1 0
0
12 Hex Display~
7 535 146 0 18 19
10 11 10 3 9 0 0 0 0 0
0 1 1 1 1 0 0 1 3
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
2 D3
-8 -38 6 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
7361 0 0
2
41149.1 0
0
12 Hex Display~
7 582 146 0 18 19
10 15 14 12 26 0 0 0 0 0
0 0 1 1 0 0 0 0 1
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
2 D2
-8 -38 6 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 512 0 0 0 0
4 DISP
4747 0 0
2
41149.1 0
0
10 2-In NAND~
219 653 409 0 3 22
0 14 12 13
0
0 0 624 512
4 7400
-7 -24 21 -16
3 ND2
-8 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
972 0 0
2
41149.1 0
0
6 JK RN~
219 1153 338 0 6 22
0 5 3 5 8 27 9
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
4 JK11
-14 -42 14 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 512 2 1 17 0
1 U
3472 0 0
2
41149.1 2
0
6 JK RN~
219 1063 338 0 6 22
0 5 10 5 8 28 3
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
4 JK10
-14 -42 14 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 512 2 2 16 0
1 U
9998 0 0
2
41149.1 0
0
6 JK RN~
219 888 338 0 6 22
0 5 12 5 8 29 11
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 JK8
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 512 2 2 9 0
1 U
3536 0 0
2
41149.1 4
0
6 JK RN~
219 974 337 0 6 22
0 5 11 5 8 30 10
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 JK9
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 512 2 1 8 0
1 U
4597 0 0
2
41149.1 1
0
6 JK RN~
219 768 338 0 6 22
0 5 14 5 13 31 12
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 JK7
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 512 2 1 6 0
1 U
3835 0 0
2
41149.1 0
0
6 JK RN~
219 697 338 0 6 22
0 32 15 5 13 33 14
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 JK6
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 512 2 1 5 0
1 U
3670 0 0
2
41149.1 0
0
6 JK RN~
219 626 338 0 6 22
0 5 16 5 13 34 15
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 JK5
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 512 2 1 4 0
1 U
5616 0 0
2
41149.1 0
0
12 Hex Display~
7 616 146 0 18 19
10 19 17 18 16 0 0 0 0 0
0 1 1 0 1 1 0 1 2
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
2 D1
-8 -38 6 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
9323 0 0
2
41149 0
0
6 JK RN~
219 217 338 0 6 22
0 5 20 5 21 35 19
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 JK1
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 512 2 2 3 0
1 U
317 0 0
2
41149 5
0
6 JK RN~
219 306 338 0 6 22
0 5 19 5 21 36 17
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 JK2
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 512 2 1 3 0
1 U
3108 0 0
2
41149 4
0
6 JK RN~
219 397 338 0 6 22
0 5 17 5 21 37 18
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 JK3
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 512 2 2 2 0
1 U
4299 0 0
2
41149 3
0
6 JK RN~
219 490 338 0 6 22
0 5 18 5 21 38 16
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 JK4
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 512 2 1 2 0
1 U
9672 0 0
2
41149 2
0
7 Pulser~
4 146 330 0 10 12
0 39 40 41 20 0 0 5 5 3
8
0
0 0 4656 0
0
3 CLK
-10 -28 11 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
7876 0 0
2
41149 1
0
10 2-In NAND~
219 246 409 0 3 22
0 17 16 21
0
0 0 624 512
4 7400
-7 -24 21 -16
3 ND1
-8 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
6369 0 0
2
41149 0
0
74
2 0 2 0 0 4096 0 6 0 0 2 3
1313 331
1296 331
1296 322
6 1 2 0 0 12416 0 5 2 0 0 5
1290 322
1296 322
1296 185
510 185
510 170
0 2 3 0 0 4096 0 0 4 47 0 3
1104 321
1104 510
988 510
0 2 4 0 0 12432 0 0 2 11 0 5
1388 322
1389 322
1389 180
504 180
504 170
1 0 5 0 0 4096 0 6 0 0 12 2
1320 322
1310 322
3 2 6 0 0 4224 0 7 3 0 0 3
936 436
897 436
897 427
0 1 7 0 0 8192 0 0 3 10 0 3
933 482
879 482
879 427
3 0 8 0 0 4096 0 3 0 0 20 2
888 382
888 374
4 0 7 0 0 4096 0 5 0 0 10 2
1266 370
1266 462
4 3 7 0 0 8320 0 6 4 0 0 5
1344 370
1344 462
933 462
933 501
937 501
6 1 4 0 0 12416 0 6 4 0 0 4
1368 322
1388 322
1388 492
988 492
0 3 5 0 0 4096 0 0 6 33 0 4
1116 274
1310 274
1310 340
1320 340
1 0 5 0 0 0 0 5 0 0 14 2
1242 322
1221 322
3 0 5 0 0 0 0 5 0 0 12 3
1242 340
1221 340
1221 274
6 2 9 0 0 12288 0 0 5 17 0 4
1187 321
1208 321
1208 331
1235 331
4 0 8 0 0 0 0 12 0 0 20 4
1063 369
1063 375
1065 375
1065 374
0 2 9 0 0 12288 0 0 7 21 0 4
1186 321
1187 321
1187 445
987 445
0 1 10 0 0 4096 0 0 7 23 0 3
1008 320
1008 427
987 427
4 0 8 0 0 0 0 14 0 0 20 2
974 368
974 374
4 4 8 0 0 8320 0 11 13 0 0 4
1153 369
1153 374
888 374
888 369
4 6 9 0 0 8320 0 8 11 0 0 5
526 170
526 190
1186 190
1186 321
1177 321
3 0 3 0 0 8320 0 8 0 0 47 4
532 170
532 196
1095 196
1095 321
2 0 10 0 0 8320 0 8 0 0 48 4
538 170
538 201
1008 201
1008 320
1 0 11 0 0 8320 0 8 0 0 49 4
544 170
544 206
921 206
921 321
0 2 12 0 0 4096 0 0 13 37 0 4
804 321
842 321
842 330
857 330
1 0 5 0 0 0 0 13 0 0 27 4
864 321
866 321
866 321
851 321
3 0 5 0 0 0 0 13 0 0 33 3
864 339
851 339
851 274
1 0 5 0 0 0 0 14 0 0 29 2
950 320
935 320
3 0 5 0 0 0 0 14 0 0 33 3
950 338
935 338
935 274
1 0 5 0 0 0 0 12 0 0 31 4
1039 321
1042 321
1042 321
1027 321
3 0 5 0 0 0 0 12 0 0 33 3
1039 339
1027 339
1027 274
1 0 5 0 0 0 0 11 0 0 33 2
1129 321
1116 321
3 0 5 0 0 12416 0 11 0 0 43 4
1129 339
1116 339
1116 274
736 274
4 0 13 0 0 4096 0 16 0 0 35 2
697 369
697 377
0 4 13 0 0 4224 0 0 15 36 0 3
626 377
768 377
768 369
4 3 13 0 0 128 0 17 10 0 0 3
626 369
626 409
628 409
0 3 12 0 0 8320 0 0 9 40 0 4
804 321
804 212
579 212
579 170
2 0 14 0 0 8320 0 9 0 0 45 4
585 170
585 218
726 218
726 321
1 0 15 0 0 12416 0 9 0 0 46 4
591 170
591 224
656 224
656 321
2 6 12 0 0 0 0 10 15 0 0 4
679 418
804 418
804 321
792 321
0 1 14 0 0 0 0 0 10 45 0 3
731 330
731 400
679 400
1 0 5 0 0 0 0 15 0 0 43 2
744 321
736 321
0 3 5 0 0 128 0 0 15 55 0 4
441 274
736 274
736 339
744 339
3 0 5 0 0 0 0 16 0 0 43 3
673 339
666 339
666 274
6 2 14 0 0 0 0 16 15 0 0 4
721 321
726 321
726 330
737 330
6 2 15 0 0 0 0 17 16 0 0 4
650 321
656 321
656 330
666 330
6 2 3 0 0 128 0 12 11 0 0 4
1087 321
1107 321
1107 330
1122 330
6 2 10 0 0 128 0 14 12 0 0 4
998 320
1021 320
1021 330
1032 330
6 2 11 0 0 128 0 13 14 0 0 4
912 321
927 321
927 329
943 329
1 0 5 0 0 0 0 17 0 0 51 2
602 321
584 321
3 0 5 0 0 0 0 17 0 0 43 3
602 339
584 339
584 274
0 2 16 0 0 8192 0 0 17 60 0 3
526 331
526 330
595 330
6 0 17 0 0 4096 0 20 0 0 57 2
330 321
347 321
0 3 18 0 0 8320 0 0 18 72 0 4
431 322
431 259
613 259
613 170
1 1 5 0 0 128 0 1 22 0 0 8
159 275
184 275
184 274
442 274
442 323
442 323
442 321
466 321
0 1 19 0 0 8320 0 0 18 71 0 4
252 321
252 253
625 253
625 170
0 2 17 0 0 8320 0 0 18 59 0 4
347 331
347 248
619 248
619 170
4 2 20 0 0 12416 0 23 19 0 0 4
176 330
174 330
174 330
186 330
2 1 17 0 0 128 0 21 24 0 0 4
366 330
347 330
347 400
272 400
0 2 16 0 0 8320 0 0 24 63 0 3
526 320
526 418
272 418
4 0 21 0 0 4096 0 19 0 0 62 2
217 369
217 379
4 3 21 0 0 8320 0 22 24 0 0 5
490 369
490 379
217 379
217 409
221 409
4 6 16 0 0 0 0 18 22 0 0 5
607 170
607 242
526 242
526 321
514 321
0 3 5 0 0 0 0 0 22 55 0 3
442 323
442 339
466 339
1 0 5 0 0 0 0 19 0 0 66 2
193 321
184 321
3 0 5 0 0 0 0 19 0 0 55 3
193 339
184 339
184 274
1 0 5 0 0 0 0 20 0 0 68 2
282 321
270 321
0 3 5 0 0 0 0 0 20 55 0 3
270 274
270 339
282 339
1 0 5 0 0 0 0 21 0 0 70 3
373 321
359 321
359 304
0 3 5 0 0 0 0 0 21 55 0 3
359 274
359 339
373 339
6 2 19 0 0 0 0 19 20 0 0 4
241 321
252 321
252 330
275 330
6 2 18 0 0 0 0 21 22 0 0 4
421 321
431 321
431 330
459 330
4 0 21 0 0 0 0 20 0 0 62 4
306 369
306 367
306 367
306 379
4 0 21 0 0 0 0 21 0 0 62 2
397 369
397 379
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 1e-06 1e-07 1e-07
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
14112 0 0 0
0
0 0 0
0
0 0 0
5 -1 10 10 10 0 10 10 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
