CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
40 10 1 100 10
176 79 1364 717
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
3 4 0.500000 0.500000
344 175 457 272
9437202 0
0
6 Title:
5 Name:
0
0
0
24
9 2-In AND~
219 195 448 0 3 22
0 2 3 18
0
0 0 624 0
6 74LS08
-21 -24 21 -16
4 U11A
-15 -25 13 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 11 0
1 U
9172 0 0
2
41143.8 0
0
10 2-In NAND~
219 259 543 0 3 22
0 5 4 2
0
0 0 624 512
4 7400
-7 -24 21 -16
4 U10D
-11 -25 17 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 10 0
1 U
7100 0 0
2
41143.8 0
0
10 2-In NAND~
219 260 488 0 3 22
0 6 7 3
0
0 0 624 512
4 7400
-7 -24 21 -16
4 U10C
-11 -25 17 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 10 0
1 U
3820 0 0
2
41143.7 0
0
10 2-In NAND~
219 231 409 0 3 22
0 13 10 11
0
0 0 624 512
4 7400
-7 -24 21 -16
4 U10B
-11 -25 17 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 10 0
1 U
7678 0 0
2
5.89581e-315 0
0
10 2-In NAND~
219 233 358 0 3 22
0 15 16 17
0
0 0 112 512
4 7400
-7 -24 21 -16
4 U10A
-11 -25 17 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 10 0
1 U
961 0 0
2
5.89581e-315 0
0
6 JK RN~
219 1104 184 0 6 22
0 9 8 9 2 23 5
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U8B
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 512 2 2 8 0
1 U
3178 0 0
2
5.89581e-315 5.26354e-315
0
6 JK RN~
219 1034 193 0 6 22
0 9 7 9 2 24 8
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U9A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 512 2 1 9 0
1 U
3409 0 0
2
5.89581e-315 0
0
12 Hex Display~
7 520 51 0 16 19
10 8 5 25 26 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP3
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 512 1 0 0 0
4 DISP
3951 0 0
2
5.89581e-315 0
0
12 Hex Display~
7 554 51 0 18 19
10 19 6 4 7 0 0 0 0 0
0 1 1 0 1 1 0 1 2
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP2
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
8885 0 0
2
5.89581e-315 0
0
6 JK RN~
219 975 202 0 6 22
0 9 4 9 18 27 7
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U7A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 512 2 1 7 0
1 U
3780 0 0
2
5.89581e-315 0
0
6 JK RN~
219 911 211 0 6 22
0 9 6 9 18 28 4
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U6B
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 512 2 2 6 0
1 U
9265 0 0
2
5.89581e-315 0
0
6 JK RN~
219 816 220 0 6 22
0 9 19 9 18 29 6
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U6A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 512 2 1 6 0
1 U
9442 0 0
2
5.89581e-315 0
0
6 JK RN~
219 741 229 0 6 22
0 9 10 9 18 30 19
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U4A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 512 2 1 4 0
1 U
9424 0 0
2
5.89581e-315 0
0
12 Hex Display~
7 596 50 0 16 19
10 20 13 10 31 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 512 1 0 0 0
4 DISP
9968 0 0
2
5.89581e-315 0
0
6 JK RN~
219 660 244 0 6 22
0 9 13 9 11 32 10
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U5A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 512 2 1 5 0
1 U
9281 0 0
2
5.89581e-315 0
0
6 JK RN~
219 579 257 0 6 22
0 9 20 9 11 33 13
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U3B
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 512 2 2 3 0
1 U
8464 0 0
2
5.89581e-315 0
0
6 JK RN~
219 511 266 0 6 22
0 9 16 9 11 34 20
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U3A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 512 2 1 3 0
1 U
7168 0 0
2
5.89581e-315 0
0
7 Pulser~
4 76 338 0 10 12
0 35 36 37 12 0 0 5 5 3
7
0
0 0 4656 0
0
2 V2
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
3171 0 0
2
5.89581e-315 0
0
2 +V
167 117 118 0 1 3
0 9
0
0 0 54256 0
3 10V
-11 -22 10 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
4139 0 0
2
5.89581e-315 0
0
12 Hex Display~
7 629 50 0 18 19
10 22 15 21 16 0 0 0 0 0
0 1 1 0 1 1 0 1 2
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
4 Sami
-15 -38 13 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
6435 0 0
2
5.89581e-315 0
0
6 JK RN~
219 439 277 0 6 22
0 9 21 9 17 38 16
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U2B
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 512 2 2 2 0
1 U
5283 0 0
2
5.89581e-315 0
0
6 JK RN~
219 372 286 0 6 22
0 9 15 9 17 39 21
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U2A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 512 2 1 2 0
1 U
6874 0 0
2
5.89581e-315 0
0
6 JK RN~
219 305 295 0 6 22
0 9 22 9 17 40 15
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U1B
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 512 2 2 1 0
1 U
5305 0 0
2
5.89581e-315 0
0
6 JK RN~
219 233 304 0 6 22
0 9 12 9 17 41 22
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U1A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 512 2 1 1 0
1 U
34 0 0
2
5.89581e-315 0
0
78
1 0 2 0 0 8192 0 1 0 0 3 4
171 439
120 439
120 529
204 529
2 3 3 0 0 12416 0 1 3 0 0 4
171 457
132 457
132 488
235 488
3 4 2 0 0 12416 0 2 6 0 0 5
234 543
204 543
204 515
1104 515
1104 215
2 2 4 0 0 4224 0 2 10 0 0 3
285 552
944 552
944 194
0 1 5 0 0 12416 0 0 2 8 0 4
1133 149
1152 149
1152 534
285 534
0 1 6 0 0 8320 0 0 3 31 0 3
862 203
862 479
286 479
2 2 7 0 0 12416 0 7 3 0 0 4
1003 185
1011 185
1011 497
286 497
2 6 5 0 0 128 0 8 6 0 0 5
523 75
523 93
1133 93
1133 167
1128 167
2 1 8 0 0 8320 0 6 8 0 0 4
1073 176
1073 99
529 99
529 75
6 2 8 0 0 0 0 7 6 0 0 2
1058 176
1073 176
3 0 9 0 0 12288 0 6 0 0 41 6
1080 185
1063 185
1063 123
940 123
940 160
941 160
0 2 10 0 0 8320 0 0 4 46 0 3
693 230
693 418
257 418
0 0 11 0 0 4096 0 0 0 58 58 5
660 379
645 379
645 378
653 378
653 379
4 2 12 0 0 4224 0 18 24 0 0 4
106 338
173 338
173 296
202 296
6 1 13 0 0 12416 0 16 4 0 0 4
603 240
625 240
625 400
257 400
0 0 14 0 0 4224 0 0 0 0 0 4
751 240
752 240
752 241
753 241
2 1 15 0 0 8192 0 22 5 0 0 3
341 278
341 349
259 349
0 2 16 0 0 8320 0 0 5 50 0 3
471 260
471 367
259 367
4 0 17 0 0 4096 0 24 0 0 20 2
233 335
233 336
4 3 17 0 0 8320 0 21 5 0 0 5
439 308
439 336
205 336
205 358
208 358
4 0 2 0 0 0 0 7 0 0 3 2
1034 224
1034 515
1 0 9 0 0 0 0 6 0 0 11 2
1080 167
1063 167
0 2 7 0 0 0 0 0 7 33 0 4
997 185
1005 185
1005 185
1003 185
1 0 9 0 0 0 0 7 0 0 25 4
1010 176
1013 176
1013 177
1002 177
3 0 9 0 0 0 0 7 0 0 11 3
1010 194
1002 194
1002 123
4 0 18 0 0 4096 0 13 0 0 29 2
741 260
741 448
4 0 18 0 0 4096 0 12 0 0 29 2
816 251
816 448
4 0 18 0 0 4096 0 11 0 0 29 2
911 242
911 448
4 3 18 0 0 8320 0 10 1 0 0 3
975 233
975 448
216 448
1 0 19 0 0 8320 0 9 0 0 44 4
563 75
563 114
770 114
770 212
2 0 6 0 0 128 0 9 0 0 43 4
557 75
557 121
862 121
862 203
3 0 4 0 0 128 0 9 0 0 42 4
551 75
551 127
935 127
935 194
4 6 7 0 0 128 0 9 10 0 0 5
545 75
545 132
997 132
997 185
999 185
1 0 9 0 0 0 0 13 0 0 35 4
717 212
721 212
721 212
706 212
3 0 9 0 0 0 0 13 0 0 41 3
717 230
706 230
706 160
1 0 9 0 0 0 0 12 0 0 37 4
792 203
794 203
794 203
779 203
3 0 9 0 0 0 0 12 0 0 41 3
792 221
779 221
779 160
1 0 9 0 0 0 0 11 0 0 39 4
887 194
895 194
895 194
880 194
3 0 9 0 0 0 0 11 0 0 41 3
887 212
880 212
880 160
1 0 9 0 0 0 0 10 0 0 41 4
951 185
956 185
956 185
941 185
0 3 9 0 0 4096 0 0 10 55 0 4
681 160
941 160
941 203
951 203
6 2 4 0 0 0 0 11 10 0 0 2
935 194
944 194
6 2 6 0 0 0 0 12 11 0 0 2
840 203
880 203
6 2 19 0 0 0 0 13 12 0 0 2
765 212
785 212
0 2 10 0 0 0 0 0 13 12 0 4
693 230
699 230
699 221
710 221
6 3 10 0 0 0 0 15 14 0 0 7
684 227
693 227
693 230
693 230
693 154
593 154
593 74
1 0 9 0 0 0 0 15 0 0 48 4
636 227
620 227
620 230
614 230
0 3 9 0 0 0 0 0 15 55 0 3
614 160
614 245
636 245
2 6 20 0 0 4096 0 16 17 0 0 6
548 249
538 249
538 251
538 251
538 249
535 249
0 2 16 0 0 0 0 0 17 63 0 4
465 260
471 260
471 258
480 258
1 0 9 0 0 0 0 17 0 0 52 4
487 249
490 249
490 250
475 250
3 0 9 0 0 0 0 17 0 0 55 3
487 267
475 267
475 160
1 0 9 0 0 0 0 16 0 0 54 4
555 240
562 240
562 240
547 240
0 3 9 0 0 0 0 0 16 55 0 3
547 160
547 258
555 258
0 0 9 0 0 4096 0 0 0 76 0 3
406 160
682 160
682 161
1 0 20 0 0 12416 0 14 0 0 49 4
605 74
605 138
538 138
538 251
2 0 13 0 0 0 0 14 0 0 61 4
599 74
599 147
605 147
605 240
3 4 11 0 0 12416 0 4 15 0 0 5
206 409
204 409
204 379
660 379
660 275
4 0 11 0 0 0 0 16 0 0 58 2
579 288
579 379
4 0 11 0 0 0 0 17 0 0 58 2
511 297
511 379
6 2 13 0 0 0 0 16 15 0 0 4
603 240
605 240
605 236
629 236
3 0 21 0 0 8320 0 20 0 0 75 4
626 74
626 173
400 173
400 269
4 6 16 0 0 0 0 20 21 0 0 5
620 74
620 198
465 198
465 260
463 260
2 0 15 0 0 8320 0 20 0 0 74 4
632 74
632 182
329 182
329 278
0 1 22 0 0 8320 0 0 20 73 0 4
257 287
257 191
638 191
638 74
0 3 9 0 0 0 0 0 21 76 0 3
406 260
406 278
415 278
1 0 9 0 0 0 0 24 0 0 68 4
209 287
211 287
211 287
196 287
3 0 9 0 0 0 0 24 0 0 76 3
209 305
196 305
196 160
1 0 9 0 0 0 0 23 0 0 70 2
281 278
266 278
0 3 9 0 0 0 0 0 23 76 0 3
266 160
266 296
281 296
1 0 9 0 0 0 0 22 0 0 72 4
348 269
354 269
354 269
337 269
0 3 9 0 0 0 0 0 22 76 0 3
337 160
337 287
348 287
6 2 22 0 0 0 0 24 23 0 0 2
257 287
274 287
6 2 15 0 0 0 0 23 22 0 0 2
329 278
341 278
6 2 21 0 0 0 0 22 21 0 0 2
396 269
408 269
1 1 9 0 0 8336 0 19 21 0 0 5
117 127
117 160
406 160
406 260
415 260
4 0 17 0 0 0 0 23 0 0 20 2
305 326
305 336
4 0 17 0 0 0 0 22 0 0 20 2
372 317
372 336
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
