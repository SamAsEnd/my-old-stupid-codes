CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
120 0 30 100 10
176 79 1364 717
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
3 4 0.500000 0.500000
344 175 457 272
42991634 0
0
6 Title:
5 Name:
0
0
0
25
9 Inverter~
13 247 525 0 2 22
0 2 5
0
0 0 624 512
6 74LS04
-21 -19 21 -11
4 U11A
-8 -20 20 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 11 0
1 U
5130 0 0
2
41141.6 0
0
10 2-In NAND~
219 245 471 0 3 22
0 4 3 6
0
0 0 624 512
4 7400
-7 -24 21 -16
4 U10C
-11 -25 17 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 10 0
1 U
391 0 0
2
41141.6 0
0
10 2-In NAND~
219 245 415 0 3 22
0 13 11 20
0
0 0 624 512
4 7400
-7 -24 21 -16
4 U10B
-11 -25 17 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 10 0
1 U
3124 0 0
2
5.89581e-315 0
0
10 2-In NAND~
219 247 358 0 3 22
0 14 15 16
0
0 0 112 512
4 7400
-7 -24 21 -16
4 U10A
-11 -25 17 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 10 0
1 U
3421 0 0
2
5.89581e-315 0
0
6 JK RN~
219 1229 166 0 6 22
0 10 2 10 5 23 9
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U7B
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 512 2 2 7 0
1 U
8157 0 0
2
5.89581e-315 5.32571e-315
0
6 JK RN~
219 1162 175 0 6 22
0 10 8 10 5 24 2
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U8A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 512 2 1 8 0
1 U
5572 0 0
2
5.89581e-315 5.30499e-315
0
6 JK RN~
219 1096 184 0 6 22
0 10 7 10 5 25 8
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U8B
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 512 2 2 8 0
1 U
8901 0 0
2
5.89581e-315 5.26354e-315
0
6 JK RN~
219 1034 193 0 6 22
0 10 3 10 5 26 7
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U9A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 512 2 1 9 0
1 U
7361 0 0
2
5.89581e-315 0
0
12 Hex Display~
7 521 51 0 18 19
10 7 8 2 9 0 0 0 0 0
0 1 1 1 1 0 0 1 3
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP3
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
4747 0 0
2
5.89581e-315 0
0
12 Hex Display~
7 554 51 0 18 19
10 17 4 18 3 0 0 0 0 0
0 1 1 1 1 0 0 1 3
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP2
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
972 0 0
2
5.89581e-315 0
0
6 JK RN~
219 970 202 0 6 22
0 10 18 10 6 27 3
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U7A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 512 2 1 7 0
1 U
3472 0 0
2
5.89581e-315 0
0
6 JK RN~
219 900 211 0 6 22
0 10 4 10 6 28 18
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U6B
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 512 2 2 6 0
1 U
9998 0 0
2
5.89581e-315 0
0
6 JK RN~
219 816 220 0 6 22
0 10 17 10 6 29 4
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U6A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 512 2 1 6 0
1 U
3536 0 0
2
5.89581e-315 0
0
6 JK RN~
219 741 229 0 6 22
0 10 11 10 6 30 17
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U4A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 512 2 1 4 0
1 U
4597 0 0
2
5.89581e-315 0
0
12 Hex Display~
7 596 51 0 18 19
10 19 13 11 31 0 0 0 0 0
0 1 1 0 1 1 0 1 2
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 512 1 0 0 0
4 DISP
3835 0 0
2
5.89581e-315 0
0
6 JK RN~
219 650 247 0 6 22
0 10 13 10 20 32 11
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U5A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 512 2 1 5 0
1 U
3670 0 0
2
5.89581e-315 0
0
6 JK RN~
219 580 257 0 6 22
0 10 19 10 20 33 13
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U3B
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 512 2 2 3 0
1 U
5616 0 0
2
5.89581e-315 0
0
6 JK RN~
219 511 268 0 6 22
0 10 15 10 20 34 19
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U3A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 512 2 1 3 0
1 U
9323 0 0
2
5.89581e-315 0
0
7 Pulser~
4 159 296 0 10 12
0 35 36 37 12 0 0 5 5 3
8
0
0 0 4656 0
0
2 V2
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
317 0 0
2
5.89581e-315 0
0
2 +V
167 196 127 0 1 3
0 10
0
0 0 54256 0
3 10V
-11 -22 10 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
3108 0 0
2
5.89581e-315 0
0
12 Hex Display~
7 629 51 0 18 19
10 22 14 21 15 0 0 0 0 0
0 1 0 1 1 1 1 1 6
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
4 Sami
-15 -38 13 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
4299 0 0
2
5.89581e-315 0
0
6 JK RN~
219 439 277 0 6 22
0 10 21 10 16 38 15
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U2B
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 512 2 2 2 0
1 U
9672 0 0
2
5.89581e-315 0
0
6 JK RN~
219 372 287 0 6 22
0 10 14 10 16 39 21
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U2A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 512 2 1 2 0
1 U
7876 0 0
2
5.89581e-315 0
0
6 JK RN~
219 305 295 0 6 22
0 10 22 10 16 40 14
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U1B
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 512 2 2 1 0
1 U
6369 0 0
2
5.89581e-315 0
0
6 JK RN~
219 233 304 0 6 22
0 10 12 10 16 41 22
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U1A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 512 2 1 1 0
1 U
9172 0 0
2
5.89581e-315 0
0
83
6 1 2 0 0 12432 0 6 1 0 0 4
1186 158
1200 158
1200 525
268 525
0 2 3 0 0 12416 0 0 2 25 0 4
997 185
1009 185
1009 480
271 480
1 0 4 0 0 4224 0 2 0 0 36 3
271 462
859 462
859 203
2 4 5 0 0 12416 0 1 5 0 0 5
232 525
205 525
205 498
1229 498
1229 197
3 4 6 0 0 12416 0 2 11 0 0 5
220 471
203 471
203 440
970 440
970 233
1 6 7 0 0 8320 0 9 8 0 0 4
530 75
530 94
1058 94
1058 176
2 0 8 0 0 8320 0 9 0 0 31 4
524 75
524 100
1126 100
1126 167
3 6 2 0 0 128 0 9 6 0 0 4
518 75
518 104
1186 104
1186 158
4 6 9 0 0 8320 0 9 5 0 0 5
512 75
512 110
1264 110
1264 149
1253 149
1 0 10 0 0 4096 0 5 0 0 30 2
1205 149
1193 149
1 0 10 0 0 0 0 6 0 0 29 2
1138 158
1132 158
0 2 11 0 0 8320 0 0 3 51 0 3
693 230
693 424
271 424
4 2 12 0 0 12416 0 19 25 0 0 4
189 296
187 296
187 296
202 296
6 1 13 0 0 12416 0 17 3 0 0 4
604 240
620 240
620 406
271 406
2 1 14 0 0 4096 0 23 4 0 0 3
341 279
341 349
273 349
0 2 15 0 0 8320 0 0 4 55 0 3
471 260
471 367
273 367
4 0 16 0 0 4096 0 25 0 0 18 2
233 335
233 336
4 3 16 0 0 8320 0 22 4 0 0 5
439 308
439 336
205 336
205 358
222 358
4 0 5 0 0 0 0 8 0 0 4 2
1034 224
1034 498
4 0 5 0 0 0 0 7 0 0 4 2
1096 215
1096 498
4 0 5 0 0 0 0 6 0 0 4 2
1162 206
1162 498
6 2 2 0 0 0 0 6 5 0 0 2
1186 158
1198 158
2 6 7 0 0 0 0 7 8 0 0 2
1065 176
1058 176
1 0 10 0 0 0 0 7 0 0 28 5
1072 167
1072 165
1071 165
1071 168
1063 168
0 2 3 0 0 0 0 0 8 38 0 4
997 185
1005 185
1005 185
1003 185
1 0 10 0 0 0 0 8 0 0 27 4
1010 176
1013 176
1013 176
1002 176
3 0 10 0 0 8192 0 8 0 0 30 3
1010 194
1002 194
1002 127
3 0 10 0 0 0 0 7 0 0 30 3
1072 185
1063 185
1063 127
3 0 10 0 0 0 0 6 0 0 30 3
1138 176
1132 176
1132 127
0 3 10 0 0 8192 0 0 5 46 0 5
936 160
936 127
1193 127
1193 167
1205 167
6 2 8 0 0 0 0 7 6 0 0 2
1120 167
1131 167
4 0 6 0 0 0 0 14 0 0 5 2
741 260
741 440
4 0 6 0 0 0 0 13 0 0 5 2
816 251
816 440
4 0 6 0 0 0 0 12 0 0 5 2
900 242
900 440
1 0 17 0 0 8320 0 10 0 0 49 4
563 75
563 114
770 114
770 212
2 0 4 0 0 0 0 10 0 0 48 4
557 75
557 121
859 121
859 203
3 0 18 0 0 8320 0 10 0 0 47 4
551 75
551 127
927 127
927 194
4 6 3 0 0 128 0 10 11 0 0 5
545 75
545 132
997 132
997 185
994 185
1 0 10 0 0 0 0 14 0 0 40 4
717 212
721 212
721 212
706 212
3 0 10 0 0 0 0 14 0 0 46 3
717 230
706 230
706 160
1 0 10 0 0 0 0 13 0 0 42 4
792 203
794 203
794 203
779 203
3 0 10 0 0 0 0 13 0 0 46 3
792 221
779 221
779 160
1 0 10 0 0 0 0 12 0 0 44 4
876 194
895 194
895 194
867 194
3 0 10 0 0 0 0 12 0 0 46 3
876 212
867 212
867 160
1 0 10 0 0 0 0 11 0 0 46 4
946 185
956 185
956 185
936 185
0 3 10 0 0 0 0 0 11 60 0 4
681 160
936 160
936 203
946 203
6 2 18 0 0 0 0 12 11 0 0 2
924 194
939 194
6 2 4 0 0 0 0 13 12 0 0 2
840 203
869 203
6 2 17 0 0 0 0 14 13 0 0 2
765 212
785 212
0 2 11 0 0 0 0 0 14 12 0 3
693 230
693 221
710 221
6 3 11 0 0 0 0 16 15 0 0 5
674 230
693 230
693 149
593 149
593 75
1 0 10 0 0 0 0 16 0 0 53 2
626 230
614 230
0 3 10 0 0 0 0 0 16 60 0 3
614 160
614 248
626 248
2 6 19 0 0 4096 0 17 18 0 0 4
549 249
538 249
538 251
535 251
0 2 15 0 0 0 0 0 18 68 0 2
465 260
480 260
1 0 10 0 0 0 0 18 0 0 57 4
487 251
490 251
490 250
475 250
3 0 10 0 0 0 0 18 0 0 60 3
487 269
475 269
475 160
1 0 10 0 0 0 0 17 0 0 59 4
556 240
562 240
562 240
547 240
0 3 10 0 0 0 0 0 17 60 0 3
547 160
547 258
556 258
0 0 10 0 0 4224 0 0 0 81 46 2
406 160
682 160
1 0 19 0 0 12416 0 15 0 0 54 4
605 75
605 138
538 138
538 251
2 0 13 0 0 0 0 15 0 0 66 4
599 75
599 143
605 143
605 240
3 4 20 0 0 12416 0 3 16 0 0 6
220 415
204 415
204 379
649 379
649 278
650 278
4 0 20 0 0 0 0 17 0 0 63 2
580 288
580 379
4 0 20 0 0 0 0 18 0 0 63 2
511 299
511 379
6 2 13 0 0 0 0 17 16 0 0 4
604 240
605 240
605 239
619 239
3 0 21 0 0 8320 0 21 0 0 80 4
626 75
626 173
400 173
400 269
4 6 15 0 0 0 0 21 22 0 0 5
620 75
620 198
465 198
465 260
463 260
2 0 14 0 0 8320 0 21 0 0 79 4
632 75
632 182
329 182
329 278
0 1 22 0 0 8320 0 0 21 78 0 4
257 287
257 191
638 191
638 75
0 3 10 0 0 0 0 0 22 81 0 3
406 260
406 278
415 278
1 0 10 0 0 0 0 25 0 0 73 4
209 287
211 287
211 287
196 287
3 0 10 0 0 0 0 25 0 0 81 3
209 305
196 305
196 160
1 0 10 0 0 0 0 24 0 0 75 2
281 278
266 278
0 3 10 0 0 0 0 0 24 81 0 3
266 160
266 296
281 296
1 0 10 0 0 0 0 23 0 0 77 4
348 270
354 270
354 269
337 269
0 3 10 0 0 0 0 0 23 81 0 3
337 160
337 288
348 288
6 2 22 0 0 0 0 25 24 0 0 2
257 287
274 287
6 2 14 0 0 0 0 24 23 0 0 3
329 278
329 279
341 279
6 2 21 0 0 0 0 23 22 0 0 4
396 270
400 270
400 269
408 269
1 1 10 0 0 128 0 20 22 0 0 5
196 136
196 160
406 160
406 260
415 260
4 0 16 0 0 0 0 24 0 0 18 2
305 326
305 336
4 0 16 0 0 0 0 23 0 0 18 2
372 318
372 336
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
