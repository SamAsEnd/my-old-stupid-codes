CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 12 100 10
177 79 1364 717
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
345 175 458 272
9437202 0
0
6 Title:
5 Name:
0
0
0
13
13 Logic Switch~
5 110 194 0 1 11
0 18
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
5.8958e-315 5.32571e-315
0
13 Logic Switch~
5 109 245 0 10 11
0 17 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
391 0 0
2
5.8958e-315 5.30499e-315
0
13 Logic Switch~
5 110 288 0 1 11
0 20
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3124 0 0
2
5.8958e-315 5.26354e-315
0
13 Logic Switch~
5 114 335 0 10 11
0 2 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3421 0 0
2
5.8958e-315 0
0
7 Pulser~
4 130 89 0 10 12
0 31 32 33 19 0 0 5 5 2
7
0
0 0 4656 0
0
5 Clock
-17 -28 18 -20
0
0
0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
8157 0 0
2
5.8958e-315 5.4086e-315
0
4 4024
219 271 179 0 9 19
0 29 30 27 25 26 28 34 35 36
0
0 0 4336 0
7 First D
-24 -60 25 -52
2 A1
-7 -70 7 -62
0
15 DVDD=14;DGND=7;
69 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o] %M
0
12 type:digital
5 DIP14
19

0 1 2 12 11 9 6 5 4 3
1 2 12 11 9 6 5 4 3 0
65 0 0 512 1 0 0 0
1 U
5572 0 0
2
5.8958e-315 5.40342e-315
0
4 4024
219 273 301 0 9 19
0 19 29 23 22 24 21 37 38 39
0
0 0 4336 0
4 4024
-14 -60 14 -52
2 A2
-7 -70 7 -62
0
15 DVDD=14;DGND=7;
69 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o %4o %5o %6o %7o %8o %9o] %M
0
12 type:digital
5 DIP14
19

0 1 2 12 11 9 6 5 4 3
1 2 12 11 9 6 5 4 3 0
65 0 0 512 1 0 0 0
1 U
8901 0 0
2
5.8958e-315 5.39824e-315
0
4 4511
219 368 206 0 20 29
0 28 26 25 27 18 17 17 10 11
12 13 14 15 16 0 0 0 0 0
2
0
0 0 4336 0
4 4511
-14 -60 14 -52
2 A3
-7 -70 7 -62
0
15 DVDD=16;DGND=8;
118 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 5 4 3 14 15
9 10 11 12 13 6 2 1 7 5
4 3 14 15 9 10 11 12 13 0
65 0 0 0 1 0 0 0
1 U
7361 0 0
2
5.8958e-315 5.39306e-315
0
4 4511
219 376 328 0 14 29
0 21 24 22 23 20 2 2 3 4
5 6 7 8 9
0
0 0 4336 0
4 4511
-14 -60 14 -52
2 A4
-7 -70 7 -62
0
15 DVDD=16;DGND=8;
118 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 6 2 1 7 5 4 3 14 15
9 10 11 12 13 6 2 1 7 5
4 3 14 15 9 10 11 12 13 0
65 0 0 0 1 0 0 0
1 U
4747 0 0
2
5.8958e-315 5.38788e-315
0
9 CC 7-Seg~
183 541 183 0 18 19
10 16 15 14 13 12 11 10 40 41
1 1 0 1 1 0 1 2 2
0
0 0 21104 0
5 REDCC
16 -41 51 -33
5 DISP1
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
972 0 0
2
5.8958e-315 5.37752e-315
0
9 CC 7-Seg~
183 594 183 0 18 19
10 9 8 7 6 5 4 3 42 43
1 1 1 1 1 1 0 2 2
0
0 0 21104 0
5 REDCC
16 -41 51 -33
5 DISP2
30 -4 65 4
0
0
32 %D %1 %2 %3 %4 %5 %6 %7 %8 %9 %S
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 0
88 0 0 512 1 0 0 0
4 DISP
3472 0 0
2
5.8958e-315 5.36716e-315
0
9 2-In AND~
219 280 347 0 3 22
0 21 22 29
0
0 0 624 180
6 74LS08
-21 -24 21 -16
3 U5A
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
9998 0 0
2
5.8958e-315 5.3568e-315
0
9 2-In AND~
219 277 224 0 3 22
0 25 26 30
0
0 0 624 180
6 74LS08
-21 -24 21 -16
3 U5B
-13 -25 8 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
3536 0 0
2
5.8958e-315 5.34643e-315
0
36
6 0 2 0 0 4096 0 9 0 0 19 2
338 337
338 342
7 8 3 0 0 8320 0 11 9 0 0 3
609 219
609 346
408 346
6 9 4 0 0 8320 0 11 9 0 0 3
603 219
603 337
408 337
5 10 5 0 0 8320 0 11 9 0 0 3
597 219
597 328
408 328
4 11 6 0 0 8320 0 11 9 0 0 3
591 219
591 319
408 319
3 12 7 0 0 8320 0 11 9 0 0 3
585 219
585 310
408 310
2 13 8 0 0 8320 0 11 9 0 0 3
579 219
579 301
408 301
1 14 9 0 0 8320 0 11 9 0 0 3
573 219
573 292
408 292
8 7 10 0 0 4224 0 8 10 0 0 5
400 224
486 224
486 255
556 255
556 219
6 9 11 0 0 16512 0 10 8 0 0 5
550 219
550 251
489 251
489 215
400 215
10 5 12 0 0 4224 0 8 10 0 0 5
400 206
493 206
493 247
544 247
544 219
11 4 13 0 0 4224 0 8 10 0 0 5
400 197
498 197
498 241
538 241
538 219
3 12 14 0 0 16512 0 10 8 0 0 5
532 219
532 236
502 236
502 188
400 188
13 2 15 0 0 4224 0 8 10 0 0 5
400 179
506 179
506 232
526 232
526 219
14 1 16 0 0 4224 0 8 10 0 0 5
400 170
511 170
511 227
520 227
520 219
0 1 17 0 0 12416 0 0 2 27 0 4
330 218
321 218
321 245
121 245
5 1 18 0 0 20608 0 8 1 0 0 6
330 206
317 206
317 241
223 241
223 194
122 194
4 1 19 0 0 8320 0 5 7 0 0 4
160 89
227 89
227 292
235 292
7 1 2 0 0 24704 0 9 4 0 0 9
338 346
338 341
332 341
332 366
331 366
331 367
222 367
222 335
126 335
5 1 20 0 0 20608 0 9 3 0 0 6
338 328
326 328
326 364
225 364
225 288
122 288
0 1 21 0 0 4224 0 0 12 26 0 3
319 292
319 356
298 356
4 2 22 0 0 8192 0 7 12 0 0 4
305 310
310 310
310 338
298 338
3 4 23 0 0 4224 0 7 9 0 0 2
305 319
344 319
4 3 22 0 0 4224 0 7 9 0 0 2
305 310
344 310
5 2 24 0 0 4224 0 7 9 0 0 2
305 301
344 301
6 1 21 0 0 0 0 7 9 0 0 2
305 292
344 292
7 6 17 0 0 0 0 8 8 0 0 2
330 224
330 215
0 1 25 0 0 4224 0 0 13 31 0 3
314 188
314 233
295 233
0 2 26 0 0 4224 0 0 13 32 0 3
308 179
308 215
295 215
3 4 27 0 0 4224 0 6 8 0 0 2
303 197
336 197
4 3 25 0 0 0 0 6 8 0 0 2
303 188
336 188
5 2 26 0 0 0 0 6 8 0 0 2
303 179
336 179
6 1 28 0 0 4224 0 6 8 0 0 2
303 170
336 170
0 2 29 0 0 4096 0 0 7 36 0 4
230 311
245 311
245 310
241 310
3 2 30 0 0 8320 0 13 6 0 0 4
250 224
236 224
236 188
239 188
3 1 29 0 0 8320 0 12 6 0 0 4
253 347
230 347
230 170
233 170
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
