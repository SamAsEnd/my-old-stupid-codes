CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 110 10
176 79 1364 747
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
3 4 0.500000 0.500000
770 79 1364 747
42991634 0
0
6 Title:
5 Name:
0
0
0
25
13 Logic Switch~
5 48 524 0 10 11
0 10 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
5130 0 0
2
41139 0
0
13 Logic Switch~
5 79 506 0 10 11
0 17 0 0 0 0 0 0 0 0
1
0
0 0 28912 0
2 5V
-9 -16 5 -8
2 V5
-11 -46 3 -38
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
391 0 0
2
41138.9 0
0
10 2-In NAND~
219 231 409 0 3 22
0 5 2 3
0
0 0 624 512
4 7400
-7 -24 21 -16
4 U10B
-11 -25 17 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 10 0
1 U
3124 0 0
2
41139 0
0
10 2-In NAND~
219 233 358 0 3 22
0 7 8 9
0
0 0 112 512
4 7400
-7 -24 21 -16
4 U10A
-11 -25 17 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 10 0
1 U
3421 0 0
2
41139 0
0
6 JK RN~
219 1229 169 0 6 22
0 14 11 14 10 24 13
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U7B
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 512 2 2 7 0
1 U
8157 0 0
2
41138.9 3
0
6 JK RN~
219 1163 179 0 6 22
0 14 12 14 10 25 11
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U8A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 512 2 1 8 0
1 U
5572 0 0
2
41138.9 2
0
6 JK RN~
219 1094 184 0 6 22
0 14 15 14 10 26 12
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U8B
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 512 2 2 8 0
1 U
8901 0 0
2
41138.9 1
0
6 JK RN~
219 1034 193 0 6 22
0 14 16 14 10 27 15
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U9A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 512 2 1 9 0
1 U
7361 0 0
2
41138.9 0
0
12 Hex Display~
7 520 51 0 18 19
10 12 11 13 15 0 0 0 0 0
0 0 1 1 0 0 0 0 1
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP3
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
4747 0 0
2
41138.9 0
0
12 Hex Display~
7 554 51 0 18 19
10 18 19 20 16 0 0 0 0 0
0 0 1 1 0 0 0 0 1
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP2
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
972 0 0
2
41138.9 0
0
6 JK RN~
219 975 202 0 6 22
0 14 20 14 17 28 16
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U7A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 512 2 1 7 0
1 U
3472 0 0
2
41138.9 0
0
6 JK RN~
219 911 211 0 6 22
0 14 19 14 17 29 20
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U6B
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 512 2 2 6 0
1 U
9998 0 0
2
41138.9 0
0
6 JK RN~
219 816 220 0 6 22
0 14 18 14 17 30 19
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U6A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 512 2 1 6 0
1 U
3536 0 0
2
41138.9 0
0
6 JK RN~
219 741 229 0 6 22
0 14 2 14 17 31 18
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U4A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 512 2 1 4 0
1 U
4597 0 0
2
41138.9 0
0
12 Hex Display~
7 596 50 0 18 19
10 21 5 2 32 0 0 0 0 0
0 1 0 1 1 0 1 1 5
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 512 0 0 0 0
4 DISP
3835 0 0
2
41138.9 0
0
6 JK RN~
219 650 247 0 6 22
0 14 5 14 3 33 2
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U5A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 512 2 1 5 0
1 U
3670 0 0
2
41138.9 0
0
6 JK RN~
219 580 257 0 6 22
0 14 21 14 3 34 5
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U3B
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 512 2 2 3 0
1 U
5616 0 0
2
41138.9 0
0
6 JK RN~
219 511 268 0 6 22
0 14 8 14 3 35 21
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U3A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 512 2 1 3 0
1 U
9323 0 0
2
41138.9 0
0
7 Pulser~
4 76 338 0 10 12
0 36 37 38 4 0 0 5 5 5
7
0
0 0 4656 0
0
2 V2
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 0 0 0 0
1 V
317 0 0
2
41138.8 0
0
2 +V
167 117 118 0 1 3
0 14
0
0 0 54256 0
3 10V
-11 -22 10 -14
2 V1
-7 -32 7 -24
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 0 0
1 V
3108 0 0
2
41138.8 0
0
12 Hex Display~
7 629 50 0 18 19
10 23 7 22 8 0 0 0 0 0
0 1 0 1 1 1 1 1 6
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
4 Sami
-15 -38 13 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
4299 0 0
2
41138.8 0
0
6 JK RN~
219 439 277 0 6 22
0 14 22 14 9 39 8
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U2B
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 512 2 2 2 0
1 U
9672 0 0
2
41138.8 0
0
6 JK RN~
219 372 287 0 6 22
0 14 7 14 9 40 22
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U2A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 512 2 1 2 0
1 U
7876 0 0
2
41138.8 0
0
6 JK RN~
219 305 295 0 6 22
0 14 23 14 9 41 7
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U1B
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 7 5 10 6 8 9 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 512 2 2 1 0
1 U
6369 0 0
2
41138.8 0
0
6 JK RN~
219 233 304 0 6 22
0 14 4 14 9 42 23
0
0 0 4720 0
6 74LS73
-22 -42 20 -34
3 U1A
-11 -42 10 -34
0
15 DVCC=4;DGND=11;
64 %D [%4bi %11bi %1i %2i %3i %4i][%4bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
0
22

0 14 1 3 2 13 12 14 1 3
2 13 12 7 5 10 6 8 9 0
0 6 0
65 0 0 512 2 1 1 0
1 U
9172 0 0
2
41138.8 0
0
82
0 2 2 0 0 8320 0 0 3 50 0 3
693 230
693 418
257 418
0 0 3 0 0 12416 0 0 0 62 0 4
649 379
645 379
645 378
653 378
4 2 4 0 0 4224 0 19 25 0 0 4
106 338
173 338
173 296
202 296
6 1 5 0 0 12416 0 17 3 0 0 4
604 240
620 240
620 400
257 400
0 0 6 0 0 4224 0 0 0 0 0 4
751 240
752 240
752 241
753 241
2 1 7 0 0 8192 0 23 4 0 0 3
341 279
341 349
259 349
0 2 8 0 0 8320 0 0 4 54 0 3
471 260
471 367
259 367
4 0 9 0 0 4096 0 25 0 0 9 2
233 335
233 336
4 3 9 0 0 8320 0 22 4 0 0 5
439 308
439 336
205 336
205 358
208 358
4 0 10 0 0 4096 0 8 0 0 13 2
1034 224
1034 524
4 0 10 0 0 4096 0 7 0 0 13 2
1094 215
1094 524
4 0 10 0 0 4096 0 6 0 0 13 2
1163 210
1163 524
1 4 10 0 0 4224 0 1 5 0 0 3
60 524
1229 524
1229 200
2 6 11 0 0 8320 0 9 6 0 0 4
523 75
523 94
1187 94
1187 162
1 0 12 0 0 8320 0 9 0 0 29 5
529 75
529 88
1117 88
1117 168
1127 168
3 6 13 0 0 8320 0 9 5 0 0 5
517 75
517 101
1254 101
1254 152
1253 152
6 2 11 0 0 0 0 6 5 0 0 4
1187 162
1197 162
1197 161
1198 161
1 0 14 0 0 4096 0 5 0 0 28 2
1205 152
1193 152
1 0 14 0 0 0 0 6 0 0 27 4
1139 162
1135 162
1135 161
1132 161
6 4 15 0 0 8320 0 8 9 0 0 4
1058 176
1058 108
511 108
511 75
2 6 15 0 0 0 0 7 8 0 0 2
1063 176
1058 176
1 0 14 0 0 0 0 7 0 0 26 4
1070 167
1071 167
1071 168
1063 168
0 2 16 0 0 4096 0 0 8 37 0 4
997 185
1005 185
1005 185
1003 185
1 0 14 0 0 0 0 8 0 0 25 4
1010 176
1013 176
1013 177
1002 177
3 0 14 0 0 8192 0 8 0 0 28 3
1010 194
1002 194
1002 127
3 0 14 0 0 0 0 7 0 0 28 3
1070 185
1063 185
1063 127
3 0 14 0 0 0 0 6 0 0 28 3
1139 180
1132 180
1132 127
0 3 14 0 0 12416 0 0 5 45 0 6
941 160
940 160
940 127
1193 127
1193 170
1205 170
6 2 12 0 0 0 0 7 6 0 0 4
1118 167
1127 167
1127 171
1132 171
4 0 17 0 0 4096 0 14 0 0 33 4
741 260
741 490
784 490
784 505
4 0 17 0 0 4096 0 13 0 0 33 4
816 251
816 490
850 490
850 505
4 0 17 0 0 4096 0 12 0 0 33 2
911 242
911 505
4 1 17 0 0 8336 0 11 2 0 0 4
975 233
975 505
91 505
91 506
1 0 18 0 0 8320 0 10 0 0 48 4
563 75
563 114
770 114
770 212
2 0 19 0 0 8320 0 10 0 0 47 4
557 75
557 121
874 121
874 203
3 0 20 0 0 8320 0 10 0 0 46 4
551 75
551 127
935 127
935 194
4 6 16 0 0 8320 0 10 11 0 0 5
545 75
545 132
997 132
997 185
999 185
1 0 14 0 0 0 0 14 0 0 39 4
717 212
721 212
721 212
706 212
3 0 14 0 0 0 0 14 0 0 45 3
717 230
706 230
706 160
1 0 14 0 0 0 0 13 0 0 41 4
792 203
794 203
794 203
779 203
3 0 14 0 0 0 0 13 0 0 45 3
792 221
779 221
779 160
1 0 14 0 0 0 0 12 0 0 43 4
887 194
895 194
895 194
880 194
3 0 14 0 0 0 0 12 0 0 45 3
887 212
880 212
880 160
1 0 14 0 0 0 0 11 0 0 45 4
951 185
956 185
956 185
941 185
0 3 14 0 0 4096 0 0 11 59 0 4
681 160
941 160
941 203
951 203
6 2 20 0 0 0 0 12 11 0 0 2
935 194
944 194
6 2 19 0 0 0 0 13 12 0 0 2
840 203
880 203
6 2 18 0 0 0 0 14 13 0 0 2
765 212
785 212
0 2 2 0 0 0 0 0 14 1 0 4
693 230
699 230
699 221
710 221
6 3 2 0 0 128 0 16 15 0 0 5
674 230
693 230
693 154
593 154
593 74
1 0 14 0 0 0 0 16 0 0 52 2
626 230
614 230
0 3 14 0 0 0 0 0 16 59 0 3
614 160
614 248
626 248
2 6 21 0 0 4096 0 17 18 0 0 4
549 249
538 249
538 251
535 251
0 2 8 0 0 0 0 0 18 67 0 2
465 260
480 260
1 0 14 0 0 0 0 18 0 0 56 4
487 251
490 251
490 250
475 250
3 0 14 0 0 0 0 18 0 0 59 3
487 269
475 269
475 160
1 0 14 0 0 0 0 17 0 0 58 4
556 240
562 240
562 240
547 240
0 3 14 0 0 0 0 0 17 59 0 3
547 160
547 258
556 258
0 0 14 0 0 4224 0 0 0 80 0 3
406 160
682 160
682 161
1 0 21 0 0 12416 0 15 0 0 53 4
605 74
605 138
538 138
538 251
2 0 5 0 0 128 0 15 0 0 65 4
599 74
599 143
605 143
605 240
3 4 3 0 0 12416 0 3 16 0 0 6
206 409
204 409
204 379
649 379
649 278
650 278
4 0 3 0 0 0 0 17 0 0 62 2
580 288
580 379
4 0 3 0 0 0 0 18 0 0 62 2
511 299
511 379
6 2 5 0 0 0 0 17 16 0 0 4
604 240
605 240
605 239
619 239
3 0 22 0 0 8320 0 21 0 0 79 4
626 74
626 173
400 173
400 269
4 6 8 0 0 128 0 21 22 0 0 5
620 74
620 198
465 198
465 260
463 260
2 0 7 0 0 8320 0 21 0 0 78 4
632 74
632 182
329 182
329 278
0 1 23 0 0 8320 0 0 21 77 0 4
257 287
257 191
638 191
638 74
0 3 14 0 0 0 0 0 22 80 0 3
406 260
406 278
415 278
1 0 14 0 0 0 0 25 0 0 72 4
209 287
211 287
211 287
196 287
3 0 14 0 0 0 0 25 0 0 80 3
209 305
196 305
196 160
1 0 14 0 0 0 0 24 0 0 74 2
281 278
266 278
0 3 14 0 0 0 0 0 24 80 0 3
266 160
266 296
281 296
1 0 14 0 0 0 0 23 0 0 76 4
348 270
354 270
354 269
337 269
0 3 14 0 0 0 0 0 23 80 0 3
337 160
337 288
348 288
6 2 23 0 0 0 0 25 24 0 0 2
257 287
274 287
6 2 7 0 0 0 0 24 23 0 0 3
329 278
329 279
341 279
6 2 22 0 0 0 0 23 22 0 0 4
396 270
400 270
400 269
408 269
1 1 14 0 0 8320 0 20 22 0 0 5
117 127
117 160
406 160
406 260
415 260
4 0 9 0 0 0 0 24 0 0 9 2
305 326
305 336
4 0 9 0 0 0 0 23 0 0 9 2
372 318
372 336
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
